`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/12/09 14:37:00
// Design Name: 
// Module Name: function_generater
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module function_generater(
    output [15:0] data,
    input [7:0] control,
    input [15:0] prescaler,
    input [15:0] compare
    );
endmodule
